module Computer12(
	input clk,
	input rst
);

endmodule
